module Counter #(parameter WIDTH = 32)(
    input[WIDTH-1:0]        hot_in[15:0],
    input[WIDTH-1:0]        cold_in[15:0],
    output[WIDTH-1:0]       out[15:0]
);

endmodule